/users/course/2023F/cs613500110003/u112062525/HW1/NangateOpenCellLibrary.lef